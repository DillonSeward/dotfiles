// https://github.com/zellij-org/zellij/blob/main/example/config.kdl
// Default Themes:
// https://zellij.dev/documentation/theme-list
theme "ayu_light"
pane_frames false
simplified_ui true
scrollback_editor "/opt/homebrew/bin/nvim"

keybinds {
     normal {
        bind "Ctrl m" {
            LaunchOrFocusPlugin "session-manager" {
                floating true
                move_to_focused_tab true
            };
            SwitchToMode "Normal"
        }        

    }
    pane {
        bind "g" {
            Run "lazygit";
            SwitchToMode "normal";
        }
    }
}
